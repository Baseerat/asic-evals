// -----------------------------------------------------------------------------
// Name : baseerat_mux_wrapper.v
// Purpose : baseerat_mux wrapper
//
// -----------------------------------------------------------------------------
// Note    : This file uses Verilog-2001.
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Module declaration
// -----------------------------------------------------------------------------
module baseerat_mux_wrapper
(
  //----------------------------------------------------------------------------
  // Clock, Clock Enables and Reset.
  //----------------------------------------------------------------------------
  clk,
  resetn,

  //----------------------------------------------------------------------------
  // Mux Interface
  //----------------------------------------------------------------------------
  din0,
  din1,
  sel,

  dout

); // baseerat_mux_wrapper


//------------------------------------------------------------------------------
// Parameters
//------------------------------------------------------------------------------
parameter DATA_WIDTH = 16; //Works with multiple of 16
parameter REG_OUT = 0;

// -----------------------------------------------------------------------------
// Signal definitions
// -----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  // Clock, Clock Enable and Reset
  //----------------------------------------------------------------------------
  input   wire                          clk;
  input   wire                          resetn;

  //----------------------------------------------------------------------------
  // Mux Interface
  //----------------------------------------------------------------------------
  //Inputs
  input                [DATA_WIDTH-1:0] din0;
  input                [DATA_WIDTH-1:0] din1;
  input                                 sel;
  //Outputs
  output               [DATA_WIDTH-1:0] dout;

  //----------------------------------------------------------------------------
  // Internal Signals
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  // Main code
  // ---------------------------------------------------------------------------
  baseerat_mux_wrapper #(
      .DATA_WIDTH (DATA_WIDTH),
      .REG_OUT    (REG_OUT)
    )
    u_baseerat_mux(
    .clk        (clk),
    .resetn     (resetn),
    .din0       (din0),
    .din1       (din1),
    .sel        (sel),
    .dout       (dout)
  );

endmodule // baseerat_mux_wrapper

// -----------------------------------------------------------------------------
// End of File
// -----------------------------------------------------------------------------
