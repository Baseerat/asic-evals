// -----------------------------------------------------------------------------
// Name : baseerat_mux.v
// Purpose : General Purpose Mux
//
// -----------------------------------------------------------------------------
// Note    : This file uses Verilog-2001.
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Module declaration
// -----------------------------------------------------------------------------
module baseerat_mux
(
  //----------------------------------------------------------------------------
  // Clock, Clock Enables and Reset.
  //----------------------------------------------------------------------------
  clk,
  resetn,

  //----------------------------------------------------------------------------
  // Mux Interface
  //----------------------------------------------------------------------------
  din0,
  din1,
  sel,

  dout

); // baseerat_mux


//------------------------------------------------------------------------------
// Parameters
//------------------------------------------------------------------------------
parameter DATA_WIDTH = 16; //Works with multiple of 16
parameter REG_OUT = 0;


localparam  DATA_WIDTH_INT = (DATA_WIDTH < 16) ? DATA_WIDTH
                                               : DATA_WIDTH/16;

// -----------------------------------------------------------------------------
// Signal definitions
// -----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  // Clock, Clock Enable and Reset
  //----------------------------------------------------------------------------
  input   wire                          clk;
  input   wire                          resetn;

  //----------------------------------------------------------------------------
  // Mux Interface
  //----------------------------------------------------------------------------
  //Inputs
  input                [DATA_WIDTH-1:0] din0;
  input                [DATA_WIDTH-1:0] din1;
  input                                 sel;
  //Outputs
  output               [DATA_WIDTH-1:0] dout;

  //----------------------------------------------------------------------------
  // Internal Signals
  //----------------------------------------------------------------------------
  wire [DATA_WIDTH-1:0] dout_nxt;
  wire [DATA_WIDTH-1:0] dout_reg;
  // -----------------------------------------------------------------------------
  // Main code
  // -----------------------------------------------------------------------------
    generate
      genvar  g;

      for (g = 0; g < DATA_WIDTH_INT; g = g + 1)
      begin : g_mux
          wire [DATA_WIDTH_INT-1:0] d_nxt;
          reg  [DATA_WIDTH_INT-1:0] d_reg;

          assign d_nxt = sel   ? din0[(g*DATA_WIDTH_INT) +: DATA_WIDTH_INT]
                               : din1[(g*DATA_WIDTH_INT) +: DATA_WIDTH_INT];

         if(REG_OUT == 1)
         begin : g_reg_out
           always @(posedge clk)
           begin : p_dout_reg
               d_reg <= d_nxt;
           end
           dout[(g*DATA_WIDTH_INT) +: DATA_WIDTH_INT] = d_reg;
         end
         else
         begin: g_comb_out
           assign dout[(g*DATA_WIDTH_INT) +: DATA_WIDTH_INT] = d_nxt;
         end

      end
    endgenerate

endmodule // baseerat_mux

// -----------------------------------------------------------------------------
// End of File
// -----------------------------------------------------------------------------
